/*
* Normalizes floating-point numbers to have valid exponents.
*/
module fpu_normalize #(
    SIGN_WIDTH = 1,
    EXPONENT_WIDTH = 11,
    SIGNIFICAND_WIDTH = 52
) (
    ports
);
    
endmodule