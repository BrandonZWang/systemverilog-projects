/*
* Controls which datapath unpacked numbers are sent to.
*/
module fpu_flow #(
    SIGN_WIDTH = 1,
    EXPONENT_WIDTH = 11,
    SIGNIFICAND_WIDTH = 52
) (
    ports
);
    
endmodule