/*
* Rounds floating-point numbers according to rounding direction.
*/
module fpu_round #(
    EXPONENT_WIDTH = 11,
    SIGNIFICAND_WIDTH = 52
) (
    ports
);
    
endmodule