/*
An FPU that conforms to the standard set forth in IEEE 754-2019.
*/
module fpu_top #(
    parameters
) (
    ports
);
     
endmodule