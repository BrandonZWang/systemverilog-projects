/*
* Performs the actual addition of floating-point significands with equal exponent.
*/
module fpu_adder_core #(
    EXPONENT_WIDTH = 11,
    SIGNIFICAND_WIDTH = 52
) (
    ports
);
    
endmodule