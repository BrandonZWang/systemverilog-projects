/*
* Rounds floating-point numbers according to rounding direction.
*/
module fpu_round #(
    SIGN_WIDTH = 1,
    EXPONENT_WIDTH = 11,
    SIGNIFICAND_WIDTH = 52
) (
    ports
);
    
endmodule