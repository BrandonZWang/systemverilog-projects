/*
* Normalizes floating-point numbers to have valid exponents.
*/
module fpu_normalize #(
    EXPONENT_WIDTH = 11,
    SIGNIFICAND_WIDTH = 52
) (
    ports
);
    
endmodule