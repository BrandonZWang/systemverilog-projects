/*
* Controls which datapath unpacked numbers are sent to.
*/
module fpu_flow #(
    EXPONENT_WIDTH = 11,
    SIGNIFICAND_WIDTH = 52
) (
    ports
);
    
endmodule