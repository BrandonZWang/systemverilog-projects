/*
---- INTRO TO FLOATING POINT NUMBERS ----
--- (a.k.a. my notes on IEE 754-2019) ---

Binary floating point number - underlying representation is binary, not decimal
Subnormal number - Special defined numbers between 0 and the minimum representable number
Exception - Raised under certain conditions. See https://en.wikipedia.org/wiki/IEEE_754#Exception_handling

*/