/*
* Repacks unpacked floating-point numbers.
*/
module fpu_pack #(
    EXPONENT_WIDTH = 11,
    SIGNIFICAND_WIDTH = 52
) (
    ports
);
    
endmodule