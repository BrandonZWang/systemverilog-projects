/*
* Repacks unpacked floating-point numbers.
*/
module fpu_pack #(
    SIGN_WIDTH = 1,
    EXPONENT_WIDTH = 11,
    SIGNIFICAND_WIDTH = 52
) (
    ports
);
    
endmodule