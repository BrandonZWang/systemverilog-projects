/*
* Unpacks floating-point numbers and proves extra info.
*/
module fpu_unpack #(
    SIGN_WIDTH = 1,
    EXPONENT_WIDTH = 11,
    SIGNIFICAND_WIDTH = 52
) (
    ports
);
    
endmodule